module url

pub struct Git {}
