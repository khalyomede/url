module url

pub struct BadlyEncodedPath {
    Error
}
