module url

pub struct Other {
    pub:
        value string
}
