module url

pub struct Http {}
