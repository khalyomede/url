module url

pub struct BadlyEncodedFragment {
    Error
}
