module url

pub struct Ftps {}
