module url

pub struct Https {}
