module url

pub struct Ssh {}
