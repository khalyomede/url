module url

// Scheme represents all possible URL schemes
pub type Scheme = Http | Https | Ftp | Ftps | Ssh | Git | File | Other
