module url

pub struct MalformedScheme {
    Error
}
