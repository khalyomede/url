module url

pub struct MissingScheme {
    Error
}
