module url

pub struct File {}
