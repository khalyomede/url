module url

pub struct TraversingAboveRoot {
    Error
}
