module url

pub struct Ftp {}
