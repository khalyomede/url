module url

pub struct MissingDomain {
    Error
}
