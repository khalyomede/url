module url

pub struct BadlyEncodedQuery {
    Error
}
